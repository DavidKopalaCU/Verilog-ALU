module seven_segment (
	output [7:0] hex
);



endmodule
